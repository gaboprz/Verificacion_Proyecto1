//================================================================================
// Módulo en el que se define la interfaz para interactuar con el "Register File", 
// además de que se define el agente, el driver y el monitor para la interacción 
// con esta interfaz
//================================================================================

// Se incluye el archivo donde están definidos los tipos de paquetes
`include "transactions.sv"



//================================================================================
// Gané la ruleta!!! atte: Amanda Hernández carnet 2020023645 :)
//================================================================================

