// Importa paquetes de UVM

import uvm_pkg::*;
`include "uvm_macros.svh"